`ifndef BIT_REP_VH
`define BIT_REP_VH

`define R2_NEG_ONE 2'sb11
`define R2_ZERO    2'sb00
`define R2_POS_ONE 2'sb01
`define R2_OTHER   2'sb10

`endif
